--- !ruby/object:Save
secret_word: gbqnl
letters: ATRZ
health: 3
