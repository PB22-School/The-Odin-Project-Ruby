--- !ruby/object:Save
secret_word: gbqnl
letters: AT
health: 5
