--- !ruby/object:Save
secret_word: erpbeq
letters: ''
health: 5
